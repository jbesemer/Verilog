
`define IpcMessageWidth  64

`define SET_MASTER_CONFIG 0x01
`define SET_PROG_DECIMATOR 0x02
`define SET_PROG_BINAVG 0x03
`define SET_PROG_BOXCAR 0x04
`define SET_BINAVG_CLR 0x05
`define SET_TRIG_SRC 0x06
`define SET_TRIG_LEVEL 0x07
`define SET_EXT_TRIG_DELAY 0x08
`define SET_EXT_TRIG_EDGE 0x09
`define SET_PRE_TRIG_INDEX 0x0A
`define SET_POST_TRIG_INDEX 0x0B
`define SET_PULSE_MASTER 0x0C
`define SET_PULSE_RST 0x0D
`define SET_GAIN 0x0E
`define SET_DATA_MODE 0x0F


`define GET_ADC_COUNTS 0x80
`define GET_IS_MASTER 0x81
`define GET_PRE_TRIG_VALUE 0x82
`define GET_POST_TRIG_VALUE 0x83
`define GET_FPGA_VERSION 0x84
